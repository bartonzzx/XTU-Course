module fa_behavioral(a,b,ci,s,co);//���ǽ�λ�ļӷ���ģ�� 
       input a,b;
       input ci;
       output  s;
       output co;
// ����������Ӵ��룬���һλȫ��������
/* Begin */

/* End */

endmodule
